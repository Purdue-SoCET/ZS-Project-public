.subckt INV A Y VDD GND
Mn Y A GND GND MODN w=10u l=0.8u m=1
Mp Y A VDD VDD MODP w=20u l=0.8u m=1
.ends INV
