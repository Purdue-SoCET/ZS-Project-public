** sch_path: /home/asicfab/a/socet59/Downloads/NAND.sch
**.subckt NAND
M3 Vout a net1 GND n1 w=20u l=0.8u m=1
M4 net1 b GND GND n1 w=20u l=0.8u m=1
Vdd VDD GND 1.8
.save i(vdd)
M1 Vout a VDD VDD p1 w=40u l=0.8u m=1
M2 Vout b VDD VDD p1 w=40u l=0.8u m=1
Vin1 a GND pulse(0 1.8 0 0.05u 0.05u 5u 10u)
.save i(vin1)
Vin3 b GND pulse(0 1.8 2.5u 0.05u 0.05u 5u 10u)
.save i(vin3)
C1 Vout GND 10f m=1
**** begin user architecture code


.model n1 nmos level=49 version=3.3.0
.model p1 pmos level=49 version=3.3.0



.tran 0.01u 30u
.save all

**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
