VERSION 5.8 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

# --------- SITE DEFINITIONS ---------
SITE CoreSite
  SIZE 1 BY 1 ;
  CLASS CORE ;
  SYMMETRY X Y ;
END CoreSite

# --------- LAYER DEFINITIONS ---------

# NWELL
LAYER NWELL
  TYPE MASTERSLICE ;
  WIDTH 5.0 ;
  SPACING 5.0 ;
END NWELL

# ACTIVE
LAYER ACTIVE
  TYPE MASTERSLICE ;
  WIDTH 0.9 ;
  SPACING 1.4 ;
END ACTIVE

# NPLUS / PPLUS SELECT
LAYER NPLUS
  TYPE MASTERSLICE ;
  WIDTH 1.4 ;
  SPACING 1.4 ;
END NPLUS

LAYER PPLUS
  TYPE MASTERSLICE ;
  WIDTH 1.4 ;
  SPACING 1.4 ;
END PPLUS

# POLY
LAYER POLY
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  WIDTH 0.8 ;
  SPACING 1.0 ;
  RESISTANCE RPERSQ 35.0 ;
END POLY

# CONTACT
LAYER CONTACT
  TYPE CUT ;
  SPACING 0.9 ;
  WIDTH 0.9 ;
END CONTACT

# METAL1
LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  WIDTH 1.1 ;
  SPACING 1.1 ;
  SPACINGTABLE PARALLELRUNLENGTH
    0 1800
  WIDTH 10.0 ;
  RESISTANCE RPERSQ 0.08 ;
END M1

# VIA1
LAYER VIA1
  TYPE CUT ;
  WIDTH 1.0 ;
  SPACING 1.0 ;
END VIA1

# METAL2
LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  WIDTH 1.2 ;
  SPACING 1.2 ;
  SPACINGTABLE PARALLELRUNLENGTH
    0 1800
  WIDTH 10.0 ;

  RESISTANCE RPERSQ 0.06 ;
END M2

# --------- VIA DEFINITIONS ---------

VIA CONTACT
  LAYER CONTACT ;
    RECT 0 0 0.9 0.9 ;
  LAYER M1 ;
    RECT -0.5 -0.5 1.4 1.4 ;
  RESISTANCE 10.0 ;
END CONTACT

VIA VIA1
  LAYER VIA1 ;
    RECT 0 0 1.0 1.0 ;
  LAYER M1 ;
    RECT -0.5 -0.5 1.5 1.5 ;
  LAYER M2 ;
    RECT -0.5 -0.5 1.5 1.5 ;
  RESISTANCE 0.5 ;
END VIA1

END LIBRARY
