** sch_path: /home/asicfab/a/socet59/Downloads/Inverter.sch
**.subckt Inverter
Vdd VDD GND 1.8
.save i(vdd)
Vin Vin GND pulse(0 1.8 0 1 1 15 30)
.save i(vin)
M1 Vout Vin VDD VDD p1 w=5u l=0.18u m=1
M2 Vout Vin GND GND n1 w=5u l=0.18u m=1
C1 Vout GND 1p m=1
**** begin user architecture code


.model n1 nmos level=49 version=3.3.0
.model p1 pmos level=49 version=3.3.0


.tran 0.5 50
.save all .print Vin Vout

**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
