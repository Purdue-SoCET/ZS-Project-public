MACRO Nand
	CLASS core ;
	FOREIGN Nand 0.000 0.000 ;
	ORIGIN 0.000 0.000 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	SIZE 21.289 BY 51.103 ;

	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.380 16.775 20.280 18.675 ;
		END
	END A

	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1;
			RECT -0.180 24.068 1.720 25.968 ;
		END
	END B

	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER M1 ;
			RECT 17.988 21.970 19.888 23.870 ;
		END
	END Y

	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M1 ;
			RECT 2.600 46.247 10.600 48.247 ;
			RECT 9.919 46.250 17.919 48.250 ;
		END
	END VDD

	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M1 ;
			RECT 2.600 1.247 10.600 3.247 ;
			RECT 9.919 1.250 17.919 3.250 ;
		END
	END VSS

	OBS
		LAYER M1 ;
			RECT 8.216 30.108 10.219 48.426 ;
			RECT 4.875 23.396 6.775 30.802 ;
			RECT 11.603 14.797 13.503 30.937 ;
			RECT 11.608 21.072 18.307 22.980 ;
			RECT 5.089 1.292 6.989 10.727 ;
		LAYER POLY1 ;
			RECT 0.096 23.421 7.882 24.553 ;
			RECT 7.084 13.182 7.884 29.383 ;
			RECT 10.479 13.273 11.279 29.779 ;
			RECT 10.591 16.362 15.183 17.227 ;
			RECT 14.211 16.363 18.803 17.228 ;
	END
END NAND

